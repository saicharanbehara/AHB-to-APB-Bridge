//definitions 

`define seq_size 10

`define ADDR_WIDTH  32
`define DATA_WIDTH  32